package shared_package;
	int error_count = 0;
    int correct_count = 0;
endpackage : shared_package